library ieee;
use ieee.std_logic_1164.all;
use work.small_8_types_and_constants.all;

entity input_port is
generic
(
	WIDTH : natural := CPU_WIDTH
);
port
(
	input : in std_logic_vector(WIDTH-1 downto 0);
	databus : out std_logic_vector(WIDTH-1 downto 0);
	enable : in std_logic
);
end input_port;

architecture bhv of input_port is
begin
	process(enable,input)
	begin
		if(enable = '0') then
			databus <= (others => 'Z');
		else
			databus <= input;
		end if;
	end process;
end bhv;

